module BCD
(
    input [7:0] DATA,
    output [7:0] LEDs
);

    assign LEDs = DATA;
    
endmodule
